`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/07/23 16:12:39
// Design Name: 
// Module Name: filter_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module filter_rom(
    input           clk,
    input           rst_n,
    input   [4:0]   aa_f,
    input   [2:0]   aa_oc,
    input   [0:0]   aa_ic,
    input           cena,
    output reg      [15:0]   qa
    );
    
    
    logic [0:24][0:6-1][0:1-1][15:0] weight    = {
16'd991,  16'd1857,  -16'd3646,  16'd3555,  -16'd6358,  -16'd12275,  
16'd3801,  -16'd3049,  -16'd2065,  -16'd1372,  -16'd7891,  -16'd7521,  
-16'd7789,  -16'd5460,  -16'd1478,  16'd2058,  -16'd11055,  16'd284,  
-16'd7664,  -16'd1503,  16'd3657,  16'd4258,  -16'd8605,  16'd3425,  
-16'd12549,  16'd4046,  16'd991,  -16'd2667,  -16'd9034,  16'd9451,  

16'd6757,  -16'd3107,  -16'd5165,  16'd8398,  -16'd712,  -16'd8824,  
16'd833,  -16'd4618,  -16'd1677,  16'd4100,  -16'd11770,  16'd2845,  
16'd3703,  16'd400,  16'd4065,  16'd5599,  -16'd7096,  16'd5207,  
-16'd4971,  16'd3849,  16'd6323,  16'd7622,  -16'd3986,  16'd8499,  
-16'd11167,  16'd9,  16'd2489,  -16'd5322,  -16'd7238,  -16'd2685,  

16'd3544,  -16'd1541,  -16'd6781,  16'd6873,  16'd1422,  -16'd3334,  
16'd10200,  16'd851,  16'd3949,  16'd3554,  16'd2978,  16'd2844,  
16'd10248,  -16'd1028,  16'd5717,  16'd5411,  16'd1671,  16'd8198,  
16'd3105,  16'd7022,  16'd7834,  16'd5995,  16'd1994,  16'd3918,  
16'd5013,  16'd4473,  -16'd2335,  16'd1274,  16'd7658,  -16'd8289,  

-16'd6942,  -16'd1513,  -16'd830,  -16'd29,  16'd10590,  16'd653,  
16'd5873,  16'd1400,  16'd2101,  16'd5218,  16'd10168,  16'd4152,  
16'd303,  16'd8975,  16'd11924,  16'd6714,  16'd7742,  16'd7072,  
16'd8499,  16'd8082,  16'd675,  16'd9646,  16'd9215,  -16'd432,  
16'd2882,  -16'd2360,  -16'd5601,  16'd9237,  16'd4977,  -16'd14323,  

-16'd6098,  16'd330,  16'd7455,  16'd27,  16'd6828,  16'd1770,  
-16'd4242,  16'd4437,  16'd5778,  -16'd7120,  16'd1863,  16'd132,  
-16'd2942,  16'd214,  16'd5341,  -16'd76,  16'd5517,  16'd4910,  
16'd4598,  16'd8200,  -16'd3331,  16'd1600,  -16'd889,  -16'd869,  
-16'd1771,  16'd5855,  -16'd5034,  16'd7883,  16'd1738,  -16'd7533
        };
    
    always_ff @(posedge clk or negedge rst_n) begin : proc_
        if(~rst_n) begin
            qa <= 0;
        end else begin
            qa <= weight[aa_f][aa_oc][aa_ic];
        end
    end
    


endmodule   